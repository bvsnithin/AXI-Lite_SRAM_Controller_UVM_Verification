

interface axilite_if ();
    
endinterface: axilite_if

class axilite_transaction extends uvm_sequence_item;

    // AXI-Lite Signals

    // Constructor
    function new ( string name = "axilite_transaction");
        super.new(name);
    endfunction: new





endclass: axilite_transaction